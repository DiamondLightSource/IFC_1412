-- Conversion of raw I2C signals into events

-- Takes into account glitches and possible race conditions

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.support.all;

entity i2c_signals is
    port (
        clk_i : in std_ulogic;

        -- Inputs from I2C bus
        scl_i : in std_ulogic;
        sda_i : in std_ulogic;

        -- Decoded events
        start_o : out std_ulogic := '0';
        stop_o : out std_ulogic := '0';
        data_valid_o : out std_ulogic := '0';
        data_bit_o : out std_ulogic
    );
end;

architecture arch of i2c_signals is
    constant DEBOUNCE_DELAY : natural := 15;
    constant DESKEW_DELAY : natural := 15;

    type state_t is (
        SCL_HIGH,           -- Normal data capturing state
        SCL_LOW,            -- Quiescent state
        SCL_DESKEW          -- Allow for delayed falling edge
    );
    signal state : state_t := SCL_HIGH;

    signal scl_in : std_ulogic;
    signal sda_in : std_ulogic;
    signal captured_sda : std_ulogic := '1';
    signal deskew_counter : natural range 0 to DESKEW_DELAY;

begin
    -- Start by debouncing both inputs.  This will eliminate any transient
    -- glitches (t_SP = 50 ns) and at the same time will ensure that the slow
    -- rising edges generated by I2C don't cause unpleasant surprises.

    debounce_scl : entity work.debounce generic map (
        DEBOUNCE_DELAY => DEBOUNCE_DELAY
    ) port map (
        clk_i => clk_i,
        signal_i => scl_i,
        signal_o => scl_in
    );

    debounce_sda : entity work.debounce generic map (
        DEBOUNCE_DELAY => DEBOUNCE_DELAY
    ) port map (
        clk_i => clk_i,
        signal_i => sda_i,
        signal_o => sda_in
    );


    process (clk_i)
        procedure emit_data is
        begin
            -- On falling edge simply emit data
            data_bit_o <= captured_sda;
            data_valid_o <= '1';
            state <= SCL_LOW;
        end;

        procedure emit_start_stop is
        begin
            if captured_sda = '1' and sda_in = '0' then
                start_o <= '1';
            elsif captured_sda = '0' and sda_in = '1' then
                stop_o <= '1';
            end if;
            captured_sda <= sda_in;
            state <= SCL_HIGH;
        end;

    begin
        if rising_edge(clk_i) then
            case state is
                when SCL_LOW =>
                    -- Wait for rising edge and capture data on rising edge
                    data_valid_o <= '0';
                    if scl_in = '1' then
                        captured_sda <= sda_in;
                        state <= SCL_HIGH;
                    end if;
                when SCL_HIGH =>
                    -- Look for falling edge of SCL or change of SDA state and
                    -- handle accordingly
                    start_o <= '0';
                    stop_o <= '0';
                    if scl_in = '0' then
                        emit_data;
                    elsif sda_in /= captured_sda then
                        -- On START/STOP we need to allow for SCL/SDA skew from
                        -- zero t_HD_DAT
                        state <= SCL_DESKEW;
                        deskew_counter <= DESKEW_DELAY;
                    end if;
                when SCL_DESKEW =>
                    if scl_in = '0' then
                        emit_data;
                    elsif deskew_counter > 0 then
                        deskew_counter <= deskew_counter - 1;
                    else
                        emit_start_stop;
                    end if;
            end case;
        end if;
    end process;
end;
